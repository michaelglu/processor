module cross_stall_controller (in_top,in_bot,stall);

input[31:0]in_top,in_bot;
output stall;



endmodule