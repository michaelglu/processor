module regfile (
    clock,
    ctrl_writeEnable_1,ctrl_writeEnable_2,
    ctrl_reset, ctrl_writeReg_1,ctrl_writeReg_2,
    ctrl_readRegA_1, ctrl_readRegB_1, data_writeReg_1,
    data_readRegA_1, data_readRegB_1,
	 ctrl_readRegA_2, ctrl_readRegB_2, data_writeReg_2,
    data_readRegA_2, data_readRegB_2,
	 
	 
	 debugR1,debugR2,debugR3,debugR4,debugR5,debugR6,debugR7,debugR8,debugR9,debugR10,debugR11,debugR12,debugR13,debugR14,debugR15,debugR16,debugR17,debugR18,debugR19,debugR20,debugR21,debugR22,debugR23,debugR24,debugR25,debugR26,debugR27,debugR28,debugR29,debugR30,debugR31
);

   input clock, ctrl_writeEnable_1,ctrl_writeEnable_2, ctrl_reset;
   input [4:0] ctrl_writeReg_1, ctrl_readRegA_1, ctrl_readRegB_1,ctrl_writeReg_2, ctrl_readRegA_2, ctrl_readRegB_2;
   input [31:0] data_writeReg_1,data_writeReg_2;
	wire clockInv;
	assign clockInv=~clock;
   output [31:0] data_readRegA_1, data_readRegB_1,data_readRegA_2, data_readRegB_2;
	
	output[31:0]debugR1,debugR2,debugR3,debugR4,debugR5,debugR6,debugR7,debugR8,debugR9,debugR10,debugR11,debugR12,debugR13,debugR14,debugR15,debugR16,debugR17,debugR18,debugR19,debugR20,debugR21,debugR22,debugR23,debugR24,debugR25,debugR26,debugR27,debugR28,debugR29,debugR30,debugR31;

   /* YOUR CODE HERE */
	wire[31:0] zero,wr_1,wr_2,we_1,we_2,rA_1,rA_2,rB_1,rB_2,r0,r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16,r17,r18,r19,r20,r21,r22,r23,r24,r25,r26,r27,r28,r29,r30,r31;
	decoder writeDecoder_1(.i(ctrl_writeReg_1),.out(wr_1));
	decoder writeDecoder_2(.i(ctrl_writeReg_2),.out(wr_2));
	
	decoder readDecoderA_1(.i(ctrl_readRegA_1),.out(rA_1));
	decoder readDecoderB_1(.i(ctrl_readRegB_1),.out(rB_1));
	decoder readDecoderA_2(.i(ctrl_readRegA_2),.out(rA_2));
	decoder readDecoderB_2(.i(ctrl_readRegB_2),.out(rB_2));
	
	and(we_1[0],wr_1[0],ctrl_writeEnable_1);
	and(we_1[1],wr_1[1],ctrl_writeEnable_1);
	and(we_1[2],wr_1[2],ctrl_writeEnable_1);
	and(we_1[3],wr_1[3],ctrl_writeEnable_1);
	and(we_1[4],wr_1[4],ctrl_writeEnable_1);
	and(we_1[5],wr_1[5],ctrl_writeEnable_1);
	and(we_1[6],wr_1[6],ctrl_writeEnable_1);
	and(we_1[7],wr_1[7],ctrl_writeEnable_1);
	and(we_1[8],wr_1[8],ctrl_writeEnable_1);
	and(we_1[9],wr_1[9],ctrl_writeEnable_1);
	and(we_1[10],wr_1[10],ctrl_writeEnable_1);
	and(we_1[11],wr_1[11],ctrl_writeEnable_1);
	and(we_1[12],wr_1[12],ctrl_writeEnable_1);
	and(we_1[13],wr_1[13],ctrl_writeEnable_1);
	and(we_1[14],wr_1[14],ctrl_writeEnable_1);
	and(we_1[15],wr_1[15],ctrl_writeEnable_1);
	and(we_1[16],wr_1[16],ctrl_writeEnable_1);
	and(we_1[17],wr_1[17],ctrl_writeEnable_1);
	and(we_1[18],wr_1[18],ctrl_writeEnable_1);
	and(we_1[19],wr_1[19],ctrl_writeEnable_1);
	and(we_1[20],wr_1[20],ctrl_writeEnable_1);
	and(we_1[21],wr_1[21],ctrl_writeEnable_1);
	and(we_1[22],wr_1[22],ctrl_writeEnable_1);
	and(we_1[23],wr_1[23],ctrl_writeEnable_1);
	and(we_1[24],wr_1[24],ctrl_writeEnable_1);
	and(we_1[25],wr_1[25],ctrl_writeEnable_1);
	and(we_1[26],wr_1[26],ctrl_writeEnable_1);
	and(we_1[27],wr_1[27],ctrl_writeEnable_1);
	and(we_1[28],wr_1[28],ctrl_writeEnable_1);
	and(we_1[29],wr_1[29],ctrl_writeEnable_1);
	and(we_1[30],wr_1[30],ctrl_writeEnable_1);
	and(we_1[31],wr_1[31],ctrl_writeEnable_1);
	
	and(we_2[0],wr_2[0],ctrl_writeEnable_2);
	and(we_2[1],wr_2[1],ctrl_writeEnable_2);
	and(we_2[2],wr_2[2],ctrl_writeEnable_2);
	and(we_2[3],wr_2[3],ctrl_writeEnable_2);
	and(we_2[4],wr_2[4],ctrl_writeEnable_2);
	and(we_2[5],wr_2[5],ctrl_writeEnable_2);
	and(we_2[6],wr_2[6],ctrl_writeEnable_2);
	and(we_2[7],wr_2[7],ctrl_writeEnable_2);
	and(we_2[8],wr_2[8],ctrl_writeEnable_2);
	and(we_2[9],wr_2[9],ctrl_writeEnable_2);
	and(we_2[10],wr_2[10],ctrl_writeEnable_2);
	and(we_2[11],wr_2[11],ctrl_writeEnable_2);
	and(we_2[12],wr_2[12],ctrl_writeEnable_2);
	and(we_2[13],wr_2[13],ctrl_writeEnable_2);
	and(we_2[14],wr_2[14],ctrl_writeEnable_2);
	and(we_2[15],wr_2[15],ctrl_writeEnable_2);
	and(we_2[16],wr_2[16],ctrl_writeEnable_2);
	and(we_2[17],wr_2[17],ctrl_writeEnable_2);
	and(we_2[18],wr_2[18],ctrl_writeEnable_2);
	and(we_2[19],wr_2[19],ctrl_writeEnable_2);
	and(we_2[20],wr_2[20],ctrl_writeEnable_2);
	and(we_2[21],wr_2[21],ctrl_writeEnable_2);
	and(we_2[22],wr_2[22],ctrl_writeEnable_2);
	and(we_2[23],wr_2[23],ctrl_writeEnable_2);
	and(we_2[24],wr_2[24],ctrl_writeEnable_2);
	and(we_2[25],wr_2[25],ctrl_writeEnable_2);
	and(we_2[26],wr_2[26],ctrl_writeEnable_2);
	and(we_2[27],wr_2[27],ctrl_writeEnable_2);
	and(we_2[28],wr_2[28],ctrl_writeEnable_2);
	and(we_2[29],wr_2[29],ctrl_writeEnable_2);
	and(we_2[30],wr_2[30],ctrl_writeEnable_2);
	and(we_2[31],wr_2[31],ctrl_writeEnable_2);
	
	
	
	assign zero[0]=1'b0;
	assign zero[1]=1'b0;
	assign zero[2]=1'b0;
	assign zero[3]=1'b0;
	assign zero[4]=1'b0;
	assign zero[5]=1'b0;
	assign zero[6]=1'b0;
	assign zero[7]=1'b0;
	assign zero[8]=1'b0;
	assign zero[9]=1'b0;
	assign zero[10]=1'b0;
	assign zero[11]=1'b0;
	assign zero[12]=1'b0;
	assign zero[13]=1'b0;
	assign zero[14]=1'b0;
	assign zero[15]=1'b0;
	assign zero[16]=1'b0;
	assign zero[17]=1'b0;
	assign zero[18]=1'b0;
	assign zero[19]=1'b0;
	assign zero[20]=1'b0;
	assign zero[21]=1'b0;
	assign zero[22]=1'b0;
	assign zero[23]=1'b0;
	assign zero[24]=1'b0;
	assign zero[25]=1'b0;
	assign zero[26]=1'b0;
	assign zero[27]=1'b0;
	assign zero[28]=1'b0;
	assign zero[29]=1'b0;
	assign zero[30]=1'b0;
	assign zero[31]=1'b0;
register r_0(.in(zero), .clk(clockInv),.we(1'b0), .reset(ctrl_reset),.out(r0));
register r_1(.in(we_1[1]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[1]|we_2[1]), .reset(ctrl_reset),.out(r1));
register r_2(.in(we_1[2]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[2]|we_2[2]), .reset(ctrl_reset),.out(r2));
register r_3(.in(we_1[3]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[3]|we_2[3]), .reset(ctrl_reset),.out(r3));
register r_4(.in(we_1[4]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[4]|we_2[4]), .reset(ctrl_reset),.out(r4));
register r_5(.in(we_1[5]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[5]|we_2[5]), .reset(ctrl_reset),.out(r5));
register r_6(.in(we_1[6]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[6]|we_2[6]), .reset(ctrl_reset),.out(r6));
register r_7(.in(we_1[7]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[7]|we_2[7]), .reset(ctrl_reset),.out(r7));
register r_8(.in(we_1[8]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[8]|we_2[8]), .reset(ctrl_reset),.out(r8));
register r_9(.in(we_1[9]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[9]|we_2[9]), .reset(ctrl_reset),.out(r9));
register r_10(.in(we_1[10]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[10]|we_2[10]), .reset(ctrl_reset),.out(r10));
register r_11(.in(we_1[11]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[11]|we_2[11]), .reset(ctrl_reset),.out(r11));
register r_12(.in(we_1[12]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[12]|we_2[12]), .reset(ctrl_reset),.out(r12));
register r_13(.in(we_1[13]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[13]|we_2[13]), .reset(ctrl_reset),.out(r13));
register r_14(.in(we_1[14]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[14]|we_2[14]), .reset(ctrl_reset),.out(r14));
register r_15(.in(we_1[15]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[15]|we_2[15]), .reset(ctrl_reset),.out(r15));
register r_16(.in(we_1[16]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[16]|we_2[16]), .reset(ctrl_reset),.out(r16));
register r_17(.in(we_1[17]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[17]|we_2[17]), .reset(ctrl_reset),.out(r17));
register r_18(.in(we_1[18]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[18]|we_2[18]), .reset(ctrl_reset),.out(r18));
register r_19(.in(we_1[19]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[19]|we_2[19]), .reset(ctrl_reset),.out(r19));
register r_20(.in(we_1[20]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[20]|we_2[20]), .reset(ctrl_reset),.out(r20));
register r_21(.in(we_1[21]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[21]|we_2[21]), .reset(ctrl_reset),.out(r21));
register r_22(.in(we_1[22]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[22]|we_2[22]), .reset(ctrl_reset),.out(r22));
register r_23(.in(we_1[23]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[23]|we_2[23]), .reset(ctrl_reset),.out(r23));
register r_24(.in(we_1[24]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[24]|we_2[24]), .reset(ctrl_reset),.out(r24));
register r_25(.in(we_1[25]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[25]|we_2[25]), .reset(ctrl_reset),.out(r25));
register r_26(.in(we_1[26]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[26]|we_2[26]), .reset(ctrl_reset),.out(r26));
register r_27(.in(we_1[27]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[27]|we_2[27]), .reset(ctrl_reset),.out(r27));
register r_28(.in(we_1[28]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[28]|we_2[28]), .reset(ctrl_reset),.out(r28));
register r_29(.in(we_1[29]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[29]|we_2[29]), .reset(ctrl_reset),.out(r29));
register r_30(.in(we_1[30]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[30]|we_2[30]), .reset(ctrl_reset),.out(r30));
register r_31(.in(we_1[31]?data_writeReg_1:data_writeReg_2), .clk(clockInv),.we(we_1[31]|we_2[31]), .reset(ctrl_reset),.out(r31));
	
tri_state_32 ta_1_0 (.in(r0), .oe(rA_1[0]), .out(data_readRegA_1));
tri_state_32 ta_1_1 (.in(r1), .oe(rA_1[1]), .out(data_readRegA_1));
tri_state_32 ta_1_2 (.in(r2), .oe(rA_1[2]), .out(data_readRegA_1));
tri_state_32 ta_1_3 (.in(r3), .oe(rA_1[3]), .out(data_readRegA_1));
tri_state_32 ta_1_4 (.in(r4), .oe(rA_1[4]), .out(data_readRegA_1));
tri_state_32 ta_1_5 (.in(r5), .oe(rA_1[5]), .out(data_readRegA_1));
tri_state_32 ta_1_6 (.in(r6), .oe(rA_1[6]), .out(data_readRegA_1));
tri_state_32 ta_1_7 (.in(r7), .oe(rA_1[7]), .out(data_readRegA_1));
tri_state_32 ta_1_8 (.in(r8), .oe(rA_1[8]), .out(data_readRegA_1));
tri_state_32 ta_1_9 (.in(r9), .oe(rA_1[9]), .out(data_readRegA_1));
tri_state_32 ta_1_10 (.in(r10), .oe(rA_1[10]), .out(data_readRegA_1));
tri_state_32 ta_1_11 (.in(r11), .oe(rA_1[11]), .out(data_readRegA_1));
tri_state_32 ta_1_12 (.in(r12), .oe(rA_1[12]), .out(data_readRegA_1));
tri_state_32 ta_1_13 (.in(r13), .oe(rA_1[13]), .out(data_readRegA_1));
tri_state_32 ta_1_14 (.in(r14), .oe(rA_1[14]), .out(data_readRegA_1));
tri_state_32 ta_1_15 (.in(r15), .oe(rA_1[15]), .out(data_readRegA_1));
tri_state_32 ta_1_16 (.in(r16), .oe(rA_1[16]), .out(data_readRegA_1));
tri_state_32 ta_1_17 (.in(r17), .oe(rA_1[17]), .out(data_readRegA_1));
tri_state_32 ta_1_18 (.in(r18), .oe(rA_1[18]), .out(data_readRegA_1));
tri_state_32 ta_1_19 (.in(r19), .oe(rA_1[19]), .out(data_readRegA_1));
tri_state_32 ta_1_20 (.in(r20), .oe(rA_1[20]), .out(data_readRegA_1));
tri_state_32 ta_1_21 (.in(r21), .oe(rA_1[21]), .out(data_readRegA_1));
tri_state_32 ta_1_22 (.in(r22), .oe(rA_1[22]), .out(data_readRegA_1));
tri_state_32 ta_1_23 (.in(r23), .oe(rA_1[23]), .out(data_readRegA_1));
tri_state_32 ta_1_24 (.in(r24), .oe(rA_1[24]), .out(data_readRegA_1));
tri_state_32 ta_1_25 (.in(r25), .oe(rA_1[25]), .out(data_readRegA_1));
tri_state_32 ta_1_26 (.in(r26), .oe(rA_1[26]), .out(data_readRegA_1));
tri_state_32 ta_1_27 (.in(r27), .oe(rA_1[27]), .out(data_readRegA_1));
tri_state_32 ta_1_28 (.in(r28), .oe(rA_1[28]), .out(data_readRegA_1));
tri_state_32 ta_1_29 (.in(r29), .oe(rA_1[29]), .out(data_readRegA_1));
tri_state_32 ta_1_30 (.in(r30), .oe(rA_1[30]), .out(data_readRegA_1));
tri_state_32 ta_1_31 (.in(r31), .oe(rA_1[31]), .out(data_readRegA_1));
	
tri_state_32 tb_1_0 (.in(r0), .oe(rB_1[0]), .out(data_readRegB_1));
tri_state_32 tb_1_1 (.in(r1), .oe(rB_1[1]), .out(data_readRegB_1));
tri_state_32 tb_1_2 (.in(r2), .oe(rB_1[2]), .out(data_readRegB_1));
tri_state_32 tb_1_3 (.in(r3), .oe(rB_1[3]), .out(data_readRegB_1));
tri_state_32 tb_1_4 (.in(r4), .oe(rB_1[4]), .out(data_readRegB_1));
tri_state_32 tb_1_5 (.in(r5), .oe(rB_1[5]), .out(data_readRegB_1));
tri_state_32 tb_1_6 (.in(r6), .oe(rB_1[6]), .out(data_readRegB_1));
tri_state_32 tb_1_7 (.in(r7), .oe(rB_1[7]), .out(data_readRegB_1));
tri_state_32 tb_1_8 (.in(r8), .oe(rB_1[8]), .out(data_readRegB_1));
tri_state_32 tb_1_9 (.in(r9), .oe(rB_1[9]), .out(data_readRegB_1));
tri_state_32 tb_1_10 (.in(r10), .oe(rB_1[10]), .out(data_readRegB_1));
tri_state_32 tb_1_11 (.in(r11), .oe(rB_1[11]), .out(data_readRegB_1));
tri_state_32 tb_1_12 (.in(r12), .oe(rB_1[12]), .out(data_readRegB_1));
tri_state_32 tb_1_13 (.in(r13), .oe(rB_1[13]), .out(data_readRegB_1));
tri_state_32 tb_1_14 (.in(r14), .oe(rB_1[14]), .out(data_readRegB_1));
tri_state_32 tb_1_15 (.in(r15), .oe(rB_1[15]), .out(data_readRegB_1));
tri_state_32 tb_1_16 (.in(r16), .oe(rB_1[16]), .out(data_readRegB_1));
tri_state_32 tb_1_17 (.in(r17), .oe(rB_1[17]), .out(data_readRegB_1));
tri_state_32 tb_1_18 (.in(r18), .oe(rB_1[18]), .out(data_readRegB_1));
tri_state_32 tb_1_19 (.in(r19), .oe(rB_1[19]), .out(data_readRegB_1));
tri_state_32 tb_1_20 (.in(r20), .oe(rB_1[20]), .out(data_readRegB_1));
tri_state_32 tb_1_21 (.in(r21), .oe(rB_1[21]), .out(data_readRegB_1));
tri_state_32 tb_1_22 (.in(r22), .oe(rB_1[22]), .out(data_readRegB_1));
tri_state_32 tb_1_23 (.in(r23), .oe(rB_1[23]), .out(data_readRegB_1));
tri_state_32 tb_1_24 (.in(r24), .oe(rB_1[24]), .out(data_readRegB_1));
tri_state_32 tb_1_25 (.in(r25), .oe(rB_1[25]), .out(data_readRegB_1));
tri_state_32 tb_1_26 (.in(r26), .oe(rB_1[26]), .out(data_readRegB_1));
tri_state_32 tb_1_27 (.in(r27), .oe(rB_1[27]), .out(data_readRegB_1));
tri_state_32 tb_1_28 (.in(r28), .oe(rB_1[28]), .out(data_readRegB_1));
tri_state_32 tb_1_29 (.in(r29), .oe(rB_1[29]), .out(data_readRegB_1));
tri_state_32 tb_1_30 (.in(r30), .oe(rB_1[30]), .out(data_readRegB_1));
tri_state_32 tb_1_31 (.in(r31), .oe(rB_1[31]), .out(data_readRegB_1));

tri_state_32 ta_2_0 (.in(r0), .oe(rA_2[0]), .out(data_readRegA_2));
tri_state_32 ta_2_1 (.in(r1), .oe(rA_2[1]), .out(data_readRegA_2));
tri_state_32 ta_2_2 (.in(r2), .oe(rA_2[2]), .out(data_readRegA_2));
tri_state_32 ta_2_3 (.in(r3), .oe(rA_2[3]), .out(data_readRegA_2));
tri_state_32 ta_2_4 (.in(r4), .oe(rA_2[4]), .out(data_readRegA_2));
tri_state_32 ta_2_5 (.in(r5), .oe(rA_2[5]), .out(data_readRegA_2));
tri_state_32 ta_2_6 (.in(r6), .oe(rA_2[6]), .out(data_readRegA_2));
tri_state_32 ta_2_7 (.in(r7), .oe(rA_2[7]), .out(data_readRegA_2));
tri_state_32 ta_2_8 (.in(r8), .oe(rA_2[8]), .out(data_readRegA_2));
tri_state_32 ta_2_9 (.in(r9), .oe(rA_2[9]), .out(data_readRegA_2));
tri_state_32 ta_2_10 (.in(r10), .oe(rA_2[10]), .out(data_readRegA_2));
tri_state_32 ta_2_11 (.in(r11), .oe(rA_2[11]), .out(data_readRegA_2));
tri_state_32 ta_2_12 (.in(r12), .oe(rA_2[12]), .out(data_readRegA_2));
tri_state_32 ta_2_13 (.in(r13), .oe(rA_2[13]), .out(data_readRegA_2));
tri_state_32 ta_2_14 (.in(r14), .oe(rA_2[14]), .out(data_readRegA_2));
tri_state_32 ta_2_15 (.in(r15), .oe(rA_2[15]), .out(data_readRegA_2));
tri_state_32 ta_2_16 (.in(r16), .oe(rA_2[16]), .out(data_readRegA_2));
tri_state_32 ta_2_17 (.in(r17), .oe(rA_2[17]), .out(data_readRegA_2));
tri_state_32 ta_2_18 (.in(r18), .oe(rA_2[18]), .out(data_readRegA_2));
tri_state_32 ta_2_19 (.in(r19), .oe(rA_2[19]), .out(data_readRegA_2));
tri_state_32 ta_2_20 (.in(r20), .oe(rA_2[20]), .out(data_readRegA_2));
tri_state_32 ta_2_21 (.in(r21), .oe(rA_2[21]), .out(data_readRegA_2));
tri_state_32 ta_2_22 (.in(r22), .oe(rA_2[22]), .out(data_readRegA_2));
tri_state_32 ta_2_23 (.in(r23), .oe(rA_2[23]), .out(data_readRegA_2));
tri_state_32 ta_2_24 (.in(r24), .oe(rA_2[24]), .out(data_readRegA_2));
tri_state_32 ta_2_25 (.in(r25), .oe(rA_2[25]), .out(data_readRegA_2));
tri_state_32 ta_2_26 (.in(r26), .oe(rA_2[26]), .out(data_readRegA_2));
tri_state_32 ta_2_27 (.in(r27), .oe(rA_2[27]), .out(data_readRegA_2));
tri_state_32 ta_2_28 (.in(r28), .oe(rA_2[28]), .out(data_readRegA_2));
tri_state_32 ta_2_29 (.in(r29), .oe(rA_2[29]), .out(data_readRegA_2));
tri_state_32 ta_2_30 (.in(r30), .oe(rA_2[30]), .out(data_readRegA_2));
tri_state_32 ta_2_31 (.in(r31), .oe(rA_2[31]), .out(data_readRegA_2));

tri_state_32 tb_2_0 (.in(r0), .oe(rB_2[0]), .out(data_readRegB_2));
tri_state_32 tb_2_1 (.in(r1), .oe(rB_2[1]), .out(data_readRegB_2));
tri_state_32 tb_2_2 (.in(r2), .oe(rB_2[2]), .out(data_readRegB_2));
tri_state_32 tb_2_3 (.in(r3), .oe(rB_2[3]), .out(data_readRegB_2));
tri_state_32 tb_2_4 (.in(r4), .oe(rB_2[4]), .out(data_readRegB_2));
tri_state_32 tb_2_5 (.in(r5), .oe(rB_2[5]), .out(data_readRegB_2));
tri_state_32 tb_2_6 (.in(r6), .oe(rB_2[6]), .out(data_readRegB_2));
tri_state_32 tb_2_7 (.in(r7), .oe(rB_2[7]), .out(data_readRegB_2));
tri_state_32 tb_2_8 (.in(r8), .oe(rB_2[8]), .out(data_readRegB_2));
tri_state_32 tb_2_9 (.in(r9), .oe(rB_2[9]), .out(data_readRegB_2));
tri_state_32 tb_2_10 (.in(r10), .oe(rB_2[10]), .out(data_readRegB_2));
tri_state_32 tb_2_11 (.in(r11), .oe(rB_2[11]), .out(data_readRegB_2));
tri_state_32 tb_2_12 (.in(r12), .oe(rB_2[12]), .out(data_readRegB_2));
tri_state_32 tb_2_13 (.in(r13), .oe(rB_2[13]), .out(data_readRegB_2));
tri_state_32 tb_2_14 (.in(r14), .oe(rB_2[14]), .out(data_readRegB_2));
tri_state_32 tb_2_15 (.in(r15), .oe(rB_2[15]), .out(data_readRegB_2));
tri_state_32 tb_2_16 (.in(r16), .oe(rB_2[16]), .out(data_readRegB_2));
tri_state_32 tb_2_17 (.in(r17), .oe(rB_2[17]), .out(data_readRegB_2));
tri_state_32 tb_2_18 (.in(r18), .oe(rB_2[18]), .out(data_readRegB_2));
tri_state_32 tb_2_19 (.in(r19), .oe(rB_2[19]), .out(data_readRegB_2));
tri_state_32 tb_2_20 (.in(r20), .oe(rB_2[20]), .out(data_readRegB_2));
tri_state_32 tb_2_21 (.in(r21), .oe(rB_2[21]), .out(data_readRegB_2));
tri_state_32 tb_2_22 (.in(r22), .oe(rB_2[22]), .out(data_readRegB_2));
tri_state_32 tb_2_23 (.in(r23), .oe(rB_2[23]), .out(data_readRegB_2));
tri_state_32 tb_2_24 (.in(r24), .oe(rB_2[24]), .out(data_readRegB_2));
tri_state_32 tb_2_25 (.in(r25), .oe(rB_2[25]), .out(data_readRegB_2));
tri_state_32 tb_2_26 (.in(r26), .oe(rB_2[26]), .out(data_readRegB_2));
tri_state_32 tb_2_27 (.in(r27), .oe(rB_2[27]), .out(data_readRegB_2));
tri_state_32 tb_2_28 (.in(r28), .oe(rB_2[28]), .out(data_readRegB_2));
tri_state_32 tb_2_29 (.in(r29), .oe(rB_2[29]), .out(data_readRegB_2));
tri_state_32 tb_2_30 (.in(r30), .oe(rB_2[30]), .out(data_readRegB_2));
tri_state_32 tb_2_31 (.in(r31), .oe(rB_2[31]), .out(data_readRegB_2));
	
	

assign debugR1=r1;
assign debugR2=r2;
assign debugR3=r3;
assign debugR4=r4;
assign debugR5=r5;
assign debugR6=r6;
assign debugR7=r7;
assign debugR8=r8;
assign debugR9=r9;
assign debugR10=r10;
assign debugR11=r11;
assign debugR12=r12;
assign debugR13=r13;
assign debugR14=r14;
assign debugR15=r15;
assign debugR16=r16;
assign debugR17=r17;
assign debugR18=r18;
assign debugR19=r19;
assign debugR20=r20;
assign debugR21=r21;
assign debugR22=r22;
assign debugR23=r23;
assign debugR24=r24;
assign debugR25=r25;
assign debugR26=r26;
assign debugR27=r27;
assign debugR28=r28;
assign debugR29=r29;
assign debugR30=r30;
assign debugR31=r31;
	
//	mux_32 ma(.select(ctrl_readRegA), .in0(r0), .in1(r1), .in2(r2), .in3(r3),.in4(r4),.in5(r5),.in6(r6),.in7(r7),.in8(r8),.in9(r9),.in10(r10),.in11(r11),.in12(r12),.in13(r13),.in14(r14),.in15(r15),.in16(r16),.in17(r17),.in18(r18),.in19(r19),.in20(r20),.in21(r21),.in22(r22),.in23(r23),.in24(r24),.in25(r25),.in26(r26),.in27(r27),.in28(r28),.in29(r29),.in30(r30),.in31(r31),.out(data_readRegA));
//	mux_32 mb(.select(ctrl_readRegB), .in0(r0), .in1(r1), .in2(r2), .in3(r3),.in4(r4),.in5(r5),.in6(r6),.in7(r7),.in8(r8),.in9(r9),.in10(r10),.in11(r11),.in12(r12),.in13(r13),.in14(r14),.in15(r15),.in16(r16),.in17(r17),.in18(r18),.in19(r19),.in20(r20),.in21(r21),.in22(r22),.in23(r23),.in24(r24),.in25(r25),.in26(r26),.in27(r27),.in28(r28),.in29(r29),.in30(r30),.in31(r31),.out(data_readRegB));

endmodule
