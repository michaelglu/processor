module predictor (shouldTakeBranch);
output shouldTakeBranch;
assign shouldTakeBranch=1'b1;

endmodule